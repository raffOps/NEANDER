library verilog;
use verilog.vl_types.all;
entity pcup_vlg_vec_tst is
end pcup_vlg_vec_tst;
