library verilog;
use verilog.vl_types.all;
entity decod4x16_vlg_check_tst is
    port(
        cinco           : in     vl_logic;
        dez             : in     vl_logic;
        dois            : in     vl_logic;
        doze            : in     vl_logic;
        nove            : in     vl_logic;
        oito            : in     vl_logic;
        onze            : in     vl_logic;
        quatorze        : in     vl_logic;
        quatro          : in     vl_logic;
        quinze          : in     vl_logic;
        seis            : in     vl_logic;
        sete            : in     vl_logic;
        tres            : in     vl_logic;
        treze           : in     vl_logic;
        um              : in     vl_logic;
        zero            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decod4x16_vlg_check_tst;
