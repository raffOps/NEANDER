library verilog;
use verilog.vl_types.all;
entity decod3x8_vlg_vec_tst is
end decod3x8_vlg_vec_tst;
