library verilog;
use verilog.vl_types.all;
entity fulladder8bits_vlg_vec_tst is
end fulladder8bits_vlg_vec_tst;
