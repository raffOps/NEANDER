library verilog;
use verilog.vl_types.all;
entity mux4x11bit_vlg_check_tst is
    port(
        outputt         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux4x11bit_vlg_check_tst;
