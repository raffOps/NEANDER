library verilog;
use verilog.vl_types.all;
entity decod3x8_vlg_check_tst is
    port(
        cinco           : in     vl_logic;
        dois            : in     vl_logic;
        quatro          : in     vl_logic;
        seis            : in     vl_logic;
        sete            : in     vl_logic;
        tres            : in     vl_logic;
        um              : in     vl_logic;
        zero            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decod3x8_vlg_check_tst;
