library verilog;
use verilog.vl_types.all;
entity pc_up_vlg_vec_tst is
end pc_up_vlg_vec_tst;
