library verilog;
use verilog.vl_types.all;
entity mux4x11bit_vlg_vec_tst is
end mux4x11bit_vlg_vec_tst;
